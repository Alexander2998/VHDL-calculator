--*****************************************************************************
--***************************  VHDL Source Code  ******************************
--*****************************************************************************
--
--  DESIGNER NAME: Alex Chen 
--
--       LAB NAME:  <lab 2 1 bit adder>
--
--      FILE NAME:  alu_and.vhd
--
-------------------------------------------------------------------------------
--
--  DESCRIPTION
--
--    This design will implement the 'and' function
--
--
-------------------------------------------------------------------------------
--
--  REVISION HISTORY
--
--  _______________________________________________________________________
-- |  DATE    | USER | Ver |  Description                                  |
-- |==========+======+=====+================================================
-- |          |      |     |
-- | 09/2/2020| XXX  | 1.0 | Created
-- |          |      |     |
--
--*****************************************************************************
--*****************************************************************************

------------------------------------------------------------------------------
-- |||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||
-- ||||                                                                   ||||
-- ||||                    COMPONENT PACKAGE                              ||||
-- ||||                                                                   ||||
-- |||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||
------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;  
use work.adder_single_bit_structural_pkg.all;

entity alu_and is 

port(input1,input2: in std_logic; 
DataOut: out std_logic);
end entity; 

architecture structure of alu_and is 
begin 
	DataOut<=(input1 and input2); 
end structure; 